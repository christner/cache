-- Created by @(#)$CDS: vhdlin version 6.1.7-64b 09/27/2016 19:46 (sjfhw304) $
-- on Sun Dec  3 17:08:40 2017


library STD;
library IEEE;

use IEEE.std_logic_1164.all;

entity jkff is port (
    J   : in  std_logic;
    K   : in  std_logic;
    Clk : in  std_logic;
    rst : in  std_logic;
    Q   : out std_logic);
end jkff;
