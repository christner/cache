-- Created by @(#)$CDS: vhdlin version 6.1.7-64b 09/27/2016 19:46 (sjfhw304) $
-- on Sun Dec  3 17:08:40 2017


architecture structural of and_4 is
begin

  output <= input4 and input3 and input2 and input1;

end structural;
