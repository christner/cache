-- Created by @(#)$CDS: vhdlin version 6.1.7-64b 09/27/2016 19:46 (sjfhw304) $
-- on Sat Dec  9 20:28:39 2017


architecture structural of or_2 is
begin

  output <= input2 or input1;

end structural;
