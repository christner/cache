-- Created by @(#)$CDS: vhdlin version 6.1.7-64b 09/27/2016 19:46 (sjfhw304) $
-- on Sun Dec  3 17:08:40 2017


library STD;
library IEEE;

use IEEE.std_logic_1164.all;

entity and_8 is port (
    input1: in  std_logic;
    input2: in  std_logic;
    input3: in  std_logic;
    input4: in  std_logic;
    input5: in  std_logic;
    input6: in  std_logic;
    input7: in  std_logic;
    input8: in  std_logic;
    output: out std_logic);
end and_8;
