-- Created by @(#)$CDS: vhdlin version 6.1.7-64b 09/27/2016 19:46 (sjfhw304) $
-- on Sun Dec  3 17:08:40 2017


architecture structural of or_4 is
begin

  output <= input4 or input3 or input2 or input1;

end structural;
